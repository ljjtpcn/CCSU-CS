LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY lpm_ram_io0 IS
PORT
(
address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
we : IN STD_LOGIC  := '1';
inclock : IN STD_LOGIC ;
outclock : IN STD_LOGIC ;
outenab : IN STD_LOGIC  := '1';
dio : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END lpm_ram_io0;


ARCHITECTURE SYN OF lpm_ram_io0 IS




COMPONENT lpm_ram_io
GENERIC (
intended_device_family : STRING;
lpm_width : NATURAL;
lpm_widthad : NATURAL;
lpm_file:STRING;
lpm_indata : STRING;
lpm_address_control : STRING;
lpm_outdata : STRING;
use_eab : STRING;
lpm_type : STRING
);
PORT (
outenab : IN STD_LOGIC ;
outclock : IN STD_LOGIC ;
address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
dio : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
inclock : IN STD_LOGIC ;
we : IN STD_LOGIC 
);
END COMPONENT;

BEGIN

lpm_ram_io_component : lpm_ram_io
GENERIC MAP (
intended_device_family => "MAX3000A",
lpm_width => 8,
lpm_widthad => 8,
lpm_file =>"initial_file.mif",
lpm_indata => "REGISTERED",
lpm_address_control => "REGISTERED",
lpm_outdata => "REGISTERED",
use_eab => "ON",
lpm_type => "LPM_RAM_IO"
)
PORT MAP (
outenab => outenab,
outclock => outclock,
address => address,
inclock => inclock,
we => we,
dio => dio
);



END SYN;
