--�����ǰ����������
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--�����ǰ������ʵ������
ENTITY H_adder IS
PORT (in_a, in_b   : IN STD_LOGIC;
      out_s, out_co: OUT STD_LOGIC);
END H_adder ;

--�����ǰ�����ṹ�������������
--ARCHITECTURE Dataflow OF H_adder IS
--BEGIN
--	out_s<= in_a XOR in_b;
--	out_co<= in_a AND in_b;
--END Dataflow;

--�����ǰ�����ṹ����Ϊ����
ARCHITECTURE Dataflow OF H_adder IS
BEGIN 
	out_s<= '1' WHEN (in_a= '0' AND in_b= '1') ELSE
	            '1' WHEN (in_a= '1' AND in_b= '0') ELSE
				'0';
	out_co<= '1' WHEN (in_a= '1' AND in_b= '1') ELSE
	            '0';
END Dataflow; 