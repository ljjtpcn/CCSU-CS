LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY fsmctrl is 
    generic(N:integer:=50000; X:integer:=10 ; Y:integer:=100); -- pin21 100Khz N for clk input freq
port(
	reset:in std_logic;--------------------------------��λreset 
	clk:in std_logic;--------------------------------ʱ���ź�
	clkcnt:out std_logic;--------------------------------ʱ���ź�
	clkfresh:out std_logic;--------------------------------ʱ���ź�
	test:out std_logic_vector(7 downto 0);--------------�����
	en_idec:out std_logic;--------------------------------ʱ���ź�
	opcode:in std_logic_vector(3 downto 0);--------------�����
	oprdata:in std_logic_vector(3 downto 0);--------------�����
	
	mcode:out std_logic_vector(21 downto 0)--------------�����
);
END fsmctrl;


Architecture RTL of fsmctrl is

TYPE State_type IS (A, B, C, D,E,F,G);  -- ����״̬
SIGNAL State : State_Type;    -- �����ź� 
SIGNAL stest: std_logic_vector(7 downto 0);--------------�����
signal ctick,clk_state,clk_fresh:std_logic;
BEGIN 

-- ����2hz clk2hz
PROCESS(clk) --����2hz�ź� tick
variable cnt1 : INTEGER RANGE 0 TO N -1; 
BEGIN 
    IF clk='1' AND clk'event THEN 
		IF cnt1=N -1 THEN 
			cnt1:=0; 
		ELSE 
			IF 	cnt1<N/2 THEN 
				ctick<='1'; 
			ELSE 
				ctick<='0';
			END IF; 
			cnt1:=cnt1+1; 
		END IF; 
	END IF; 
end process; 

PROCESS(ctick) --����1hz�ź� clk_state
BEGIN 
   IF (reset ='0') THEN
       clk_state<='1';
	ELSIF ctick='1' AND ctick'event THEN 
		clk_state<=not clk_state; 
	END IF; 
end process; 


-- ����10khz clk10khz
PROCESS(clk) --����10Khz�ź� 
variable cnt1 : INTEGER RANGE 0 TO X -1; 
BEGIN 
	IF rising_edge(clk) THEN 
		IF cnt1=X -1 THEN 
			cnt1:=0; 
		ELSE 
			IF 	cnt1<X/2 THEN 
				clk_fresh<='1'; 
			ELSE 
				clk_fresh<='0'; 
			END IF; 
			cnt1:=cnt1+1; 
		END IF; 
	END IF; 
end process; 

  PROCESS (clk_state, reset,opcode) 
  CONSTANT LDA:std_logic_vector(3 downto 0):="0000" ;-- LDA:=0010
  CONSTANT ADD:std_logic_vector(3 downto 0):="0111" ; -- ADD:=1100 
  CONSTANT YAND:std_logic_vector(3 downto 0):="1110" ; -- YAND:=1110
  CONSTANT JMP:std_logic_vector(3 downto 0):="0101" ; -- JMP:=0001
  CONSTANT SUB:std_logic_vector(3 downto 0):="0011" ;-- sub:=0110
  CONSTANT com:std_logic_vector(3 downto 0):="0110" ; -- INC :=0111
  CONSTANT STA:std_logic_vector(3 downto 0):="1000" ; -- INC :=0111
  

  variable vmcode: std_logic_vector(21 downto 0);
  
  variable ven_idec: std_logic;
  BEGIN  
--21sw-20r4-19r5-18alu-17pc|16r1-15r2-14r4-13r5-12ar|11m-10cn-9s38s27s16s0|5pcclr-4pcld-3pcen|2memen-1mw-0mr
--   x_busLD...������P Cmem 
--      a            c
--   srrlprrrra csssslleewr
--   w45uc1245rmn3210rdnnrd
--  "1111100000000000100100"
--  "1111100001000000100101"
    If (reset = '0') THEN            -- ��λreset����λ״̬ΪA
		State <= A;
		vmcode :="1111100000000000100100";--  
		ven_idec:='0';--��������
		stest <="00000000";
    ELSIF rising_edge(clk_state) THEN   
		ven_idec:='0';
		vmcode :="1111100000000000100100";
		CASE State IS
			WHEN A => 
				vmcode :="1111000001000000111100";--  PC=>AR,PC++
				stest <="00000001";
				State <= B; 

			WHEN B => 
				vmcode :="1111100100000000100101";--  M=>r4(r4ָ��Ĵ���)
				ven_idec:='1';     --����������
				stest <="00000010";
				State <= C; 
			WHEN C => 
				CASE opcode IS
				when  LDA => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				
				when  STA => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				when  ADD => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				when  JMP => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				when  SUB => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				when  COM => vmcode :="1111000001000000111100";--  PC=>AR,PC++
				WHEN others =>NULL;
				END CASE;
				stest <="00000011";
				State <= D; 
			WHEN D => 
				CASE opcode IS
				when LDA => vmcode :="1111100001000000100101";--  M=>ar
				when COM => vmcode :="1111100001000000100101";--  M=>ar
				when ADD => vmcode :="1111100001000000100101";--  M=>ar
				when SUB => vmcode :="1111100001000000100101";--  M=>ar
				when JMP => vmcode :="1111100000000000101101";--  M=>PC
				when STA => vmcode :="1111100001000000100101";--  M=>ar
				
				WHEN others =>NULL;
				END CASE;
				stest <="00000100";
				State <= E; 
		WHEN E => 
				CASE opcode IS
				 WHEN LDA => vmcode :="1111100010000000100101";
				 WHEN COM => vmcode :="1111110000000000100101";
				 WHEN ADD => vmcode :="1111101000000000100101";
				 WHEN SUB => vmcode :="1111101000000000100101";
				 WHEN STA => vmcode :="1101100000000000100110";
				WHEN others =>NULL;
				END CASE;
				stest <="00000101";
				State <= F; 
		
			WHEN F => 
				CASE opcode IS
				 
				 WHEN ADD => vmcode :="1101110000000000100100";
				 WHEN SUB => vmcode :="1101
				 ..110000000000100100";
				WHE9++9+N others =>NULL;
				END CASE;
				stest <="00000110";
				State <= G; 
			
			WHEN G=> 
				CASE opcode IS
				 WHEN ADD => vmcode :="1110100010011001100100";
				 WHEN SUB => vmcode :="1110100010000110100100";
				 WHEN COM => vmcode :="1110100010100000100100";
				WHEN others =>NULL;
				END CASE;
				stest <="00000111";
				State <= A;
			
			WHEN others =>NULL;
		END CASE; 
    END IF; 
    mcode <=vmcode;
    en_idec <=ven_idec;
END PROCESS;
test <=stest;
clkcnt <= ctick;
clkfresh<=clk_fresh;
END rtl;

 
