LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--LIBRARY work;
LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY datapath IS
port(
	reset:in std_logic; --ʱ�� 
	clk:in std_logic; --ʱ�� 
	k:in std_logic_vector(7 downto 0);--����ʾ���ƣ�abcdefg�� 
	seg:out std_logic_vector(7 downto 0);--����ʾ���ƣ�abcdefg�� 
	y:out std_logic_vector(7 downto 0); --����ܵ�ַѡ����� 
	dout:inout std_logic_vector(7 downto 0) --����ܵ�ַѡ����� 
);
END datapath;

ARCHITECTURE Structural OF datapath IS

--ATTRIBUTE black_box : BOOLEAN;
--nATTRIBUTE noopt : BOOLEAN;

--COMPONENT lpm_ram_io_0
--	PORT(memenab : IN STD_LOGIC;
--		 inclock : IN STD_LOGIC;
--		 we : IN STD_LOGIC;
--		 outenab : IN STD_LOGIC;
--		 address : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
--);
--END COMPONENT;
--ATTRIBUTE black_box OF lpm_ram_io_0: COMPONENT IS true;
--ATTRIBUTE noopt OF lpm_ram_io_0: COMPONENT IS true;

COMPONENT idec IS
PORT(  clk,reset,en_idec:IN STD_LOGIC;
	   oprdata :out    STD_LOGIC_VECTOR(3 DOWNTO 0);
	   opcode  :OUT   STD_LOGIC_VECTOR(3 DOWNTO 0);
	   instruction      :INOUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
END COMPONENT;

COMPONENT lpm_ram_io0 IS
PORT
(
address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
we : IN STD_LOGIC  := '1';
inclock : IN STD_LOGIC ;
outclock : IN STD_LOGIC ;
outenab : IN STD_LOGIC  := '1';
dio : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END COMPONENT;

COMPONENT exp_r_alu is
port(	clk,reset                    :IN STD_LOGIC;
		sw_bus,r4_bus,r5_bus,alu_bus,memen :IN STD_LOGIC;
		lddr1,lddr2,ldr4,ldr5        :IN STD_LOGIC;
		m,cn                         :IN STD_LOGIC;
		s                            :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		k                            :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		d                            :INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
 );
END COMPONENT;

 
COMPONENT sw_pc_ar IS
PORT(  clk,pcclr,pcld,pcen,reset:IN STD_LOGIC;
	   sw_bus,pc_bus,ldar,memen     :IN STD_LOGIC;
	   inputd :IN    STD_LOGIC_VECTOR(7 DOWNTO 0);
	   arout  :OUT   STD_LOGIC_VECTOR(7 DOWNTO 0);
	   d      :INOUT STD_LOGIC_VECTOR(7 DOWNTO 0) 
);
END COMPONENT;



COMPONENT display is
port(
	clk:in std_logic;--------------------------------ʱ���ź�
	in84:in std_logic_vector(7 downto 0);--------------�����
	in83:in std_logic_vector(7 downto 0);--------------�����
	in82:in std_logic_vector(7 downto 0);--------------�����
	in81:in std_logic_vector(7 downto 0);--------------�����
	seg:out std_logic_vector(7 downto 0);--------------�����
	sel:out std_logic_vector(7 downto 0) -------------��λ
);
END COMPONENT;


COMPONENT fsmctrl is
port(
	reset:in std_logic;--------------------------------ʱ���ź�
	clk:in std_logic;--------------------------------ʱ���ź�
	clkcnt:out std_logic;--------------------------------ʱ���ź�
	clkfresh:out std_logic;--------------------------------ʱ���ź�
	test:out std_logic_vector(7 downto 0);
	en_idec:out std_logic;--------------------------------ʱ���ź�
	opcode:in std_logic_vector(3 downto 0);--------------�����
	oprdata:in std_logic_vector(3 downto 0);--------------�����
		
	mcode:out std_logic_vector(21 downto 0)
);
END COMPONENT;

--21bus16ld11op5pc2m
--21sw-20r4-19r5-18alu-17pc|16r1-15r2-14r4-13r5-12ar|11m-10cn-9s38s27s16s0|5pcclr-4pcld-3pcen|2memen-1mw-0mr
SIGNAL smcode: std_logic_vector(21 downto 0); 
SIGNAL clkcnt,clkread: std_logic; 
SIGNAL clkfresh: std_logic; 
SIGNAL sar: std_logic_vector(7 downto 0); 
SIGNAL sdbus: std_logic_vector(7 downto 0); 
SIGNAL smibus: std_logic_vector(7 downto 0); 
SIGNAL test: std_logic_vector(7 downto 0); 
SIGNAL s_opcode,s_oprdata: std_logic_vector(3 downto 0); 
SIGNAL s_enidec:STD_LOGIC; 

SIGNAL clkon:STD_LOGIC; 
begin

PROCESS(clkcnt) --
BEGIN 
    IF (reset ='0') THEN
       clkon<='1';
	ELSIF clkcnt='1' AND clkcnt'event THEN 
		clkon<=not clkon; 
	END IF; 
end process; 

PROCESS(clkcnt,clkon) --
BEGIN 
    IF (reset ='0') THEN
       clkread<='0';
	ELSIF clkcnt='0' AND clkcnt'event THEN 
		--if clkon='0' then
		   clkread<=not clkread; 
		--end if;
	END IF; 
end process; 


U0: fsmctrl PORT MAP (  
	reset => reset,
	   clk   =>clk,
       clkcnt => clkcnt,
       clkfresh => clkfresh,
       test =>test,
       en_idec=>s_enidec,
       opcode=>s_opcode,
       oprdata=>s_oprdata,
       mcode  => smcode
);

U1: sw_pc_ar PORT MAP (
       clk =>clkcnt,
       reset =>reset,
        memen =>smcode( 0),
       pcclr =>smcode( 5) ,
       pcld=>smcode( 4),
       pcen=>smcode( 3),
	   sw_bus=>smcode( 21),
	   pc_bus=>smcode( 17),
	   ldar=>smcode( 12),
	   inputd =>k,
	   arout =>sar,
	   d=>sdbus 
);

U_idec: idec PORT MAP (
       clk =>clkcnt,
       reset=>reset,
       en_idec=>s_enidec,
	   oprdata=>s_oprdata,
	   opcode=>s_opcode,
	   instruction=>sdbus 
);


U2: lpm_ram_io0 PORT MAP(
address =>sar,
we => smcode( 1),--and clkon
inclock  =>   clkcnt,
outclock  =>  clkcnt ,
outenab =>  smcode( 0) ,
dio =>sdbus
);


U3: exp_r_alu PORT MAP (
	    clk   =>clkcnt,
	    reset =>reset,
	    memen =>smcode( 0),
		sw_bus=>smcode( 21),
		r4_bus=>smcode( 20),
		r5_bus=>smcode( 19),
		alu_bus =>smcode( 18),
		lddr1 =>smcode( 16),
		lddr2=>smcode( 15),
		ldr4=>smcode( 14),
		ldr5  =>smcode( 13),
		m =>smcode( 11)	,
		cn   =>smcode(10),
		s   =>smcode(9 downto 6),
		k   =>k,
		d  =>sdbus
);


U4: display PORT MAP (
	clk  => clkfresh,
	in84 => test,
	in83 => sar,
	in82 => "00000000",
	in81 => sdbus,
	seg  => seg,
	sel  => y
);


end Structural;